//# 3 inputs
//# 6 outputs
//# 21 D-type flipflops
//# 59 inverters
//# 99 gates (11 ANDs + 30 NANDs + 24 ORs + 34 NORs)

module dff (CK,Q,D);
input CK,D;
output Q;
reg Q;
always @ (posedge CK)
  Q <= D;
endmodule

module s382(CK,G200,G201,G301,G302,G303,G304,G202,G305,G306);
input CK,G201,G202,G200;
output G301,G302,G303,G306,G304,G305;

  wire G0,G1,G2,G3,G4,G5,
   G6,G7,G8,G9,G10,G11,G12,G13,
   G14,G15,G16,G17,G18,G19,G20,G21,
    G22,G23,G24,G25,G26,G27,G28,G29,G30,G31,
    G32,G33,G34,G35,G36,G37,G38,G39,G40,G41,
   G42,G43,G44,G45,G46,G47,G48,
    G49,G50,G51,G52,G53,G54,G55,G56,G57,G58,G59,
    G60,G61,G62,G63,G64,G65,G66,
    G67,G68,G69,G70,
    G71,G72,G73,G74,G75,G76,G77,
    G78,G79,G80,G81,
  G82,G83,G84,G85,G86,G87,G88,G89,
  G90,G91,G92,G93,G94,G95,G96,
   G97,G98,G99,G100,G101,G102,
    G103,G104,G105,G106,
    G107,G108,G109,G110,G111,G112,
    G113,G114,G115,G116,
    G117,G118,G119,G120,
    G121,G122,G123,G124,
    G125,G126,G127,G128,G129,G130,
    G131,G132,G133,G134,G135,G136,
   G137,G138,G139,G140,G141,G142,
    G143,G144,G145,G146,G147,G148,
    G149,G150,G151,G152,G153,G154,
    G155,G156,G157,G158,G159,G160,G161,
    G162,G163,G164,G165,G166,G167,G168,G169,
    G170,G171,G172;
  wire SPL0_OUT1, SPL0_OUT2, SPL1_OUT1, SPL1_OUT2, SPL2_OUT1, SPL2_OUT2,
  SPL3_OUT1, SPL3_OUT2, SPL4_OUT1, SPL4_OUT2, SPL5_OUT1, SPL5_OUT2,
  SPL6_OUT1, SPL6_OUT2, SPL7_OUT1, SPL7_OUT2, SPL8_OUT1, SPL8_OUT2,
  SPL9_OUT1, SPL9_OUT2, SPL10_OUT1, SPL10_OUT2, SPL11_OUT1, SPL11_OUT2,
  SPL12_OUT1, SPL12_OUT2, SPL13_OUT1, SPL13_OUT2, SPL14_OUT1, SPL14_OUT2;

  spl SPL0(SPL0_OUT1, SPL0_OUT2, G0);// first level split of G0
  spl SPL1(SPL1_OUT1, SPL1_OUT2, SPL0_OUT2); //second level split of G0
  spl SPL2(SPL2_OUT1, SPL2_OUT2, G2); // cc
  spl SPL3(SPL3_OUT1, SPL3_OUT2, SPL2_OUT1); // second level split out1 of G2
  spl SPL4(SPL4_OUT1, SPL4_OUT2, SPL2_OUT2); // second level split out2 of G2
  spl SPL5(SPL5_OUT1, SPL5_OUT2, G9); // first level split of G9
  spl SPL6(SPL6_OUT1, SPL6_OUT2, --); // 
  spl SPL7(SPL7_OUT1, SPL7_OUT2, --); // 
  spl SPL8(SPL8_OUT1, SPL8_OUT2, --); // first level split of 
  spl SPL9(SPL9_OUT1, SPL9_OUT2, --); // first level split of 
  spl SPL10(SPL10_OUT1, SPL10_OUT2, --); // first level split of 
  spl SPL11(SPL11_OUT1, SPL11_OUT2,--); 

  
  

  dff DFF_0(CK,G0,G1);
  dff DFF_1(CK,G2,G3);
  dff DFF_2(CK,G4,G5);
  dff DFF_3(CK,G6,G7);
  dff DFF_4(CK,G8,SPL5_OUT1);
  dff DFF_5(CK,G10,G11);
  dff DFF_6(CK,G12,G13);
  dff DFF_7(CK,G14,G15);
  dff DFF_8(CK,G16,G17);
  dff DFF_9(CK,G18,G19);
  dff DFF_10(CK,G20,G21);
  dff DFF_11(CK,G22,G23);
  dff DFF_12(CK,G24,G25);
  dff DFF_13(CK,G26,G27);
  dff DFF_14(CK,G28,G29);
  dff DFF_15(CK,G30,G31);
  dff DFF_16(CK,G32,G33);
  dff DFF_17(CK,G34,G35);
  dff DFF_18(CK,G36,G37);
  dff DFF_19(CK,G38,G39);
  dff DFF_20(CK,G40,G41);
  not NOT_0(G42,SPL0_OUT1);
  not NOT_1(G43,SPL3_OUT1);
  not NOT_2(G44,G6);
  not NOT_3(G45,G8);
  not NOT_4(G46,G18);
  not NOT_5(G47,G20);
  not NOT_6(G48,G22);
  not NOT_7(G49,G24);
  not NOT_8(G50,G26);
  not NOT_9(G51,G28);
  not NOT_10(G52,G30);
  not NOT_11(G53,G32);
  not NOT_12(G54,G34);
  not NOT_13(G55,G36);
  not NOT_14(G56,G38);
  not NOT_15(G57,G40);
  not NOT_16(G58,G201);
  not NOT_17(G59,G200);
  not NOT_18(G60,SPL3_OUT2);
  not NOT_19(G61,G202);
  not NOT_20(G62,G24);
  not NOT_21(G63,G22);
  not NOT_22(G64,G20);
  not NOT_23(G65,G18);
  not NOT_24(G66,G40);
  not NOT_25(G67,G14);
  not NOT_26(G68,G12);
  not NOT_27(G69,G16);
  not NOT_28(G70,G10);
  not NOT_29(G71,G4);
  not NOT_30(G72,G58);
  not NOT_31(G73,G59);
  not NOT_32(G74,G61);
  not NOT_33(G75,G66);
  not NOT_34(G76,G57);
  not NOT_35(G301,G67);
  not NOT_36(G302,G68);
  not NOT_37(G303,G70);
  not NOT_38(G306,G71);
  not NOT_39(G77,G45);
  not NOT_40(G78,G44);
  not NOT_41(G79,G72);
  not NOT_42(G80,G73);
  not NOT_43(G81,G73);
  not NOT_44(G82,G73);
  not NOT_45(G83,G74);
  not NOT_46(G304,G77);
  not NOT_47(G305,G78);
  not NOT_48(G84,G85);
  not NOT_49(G86,G87);
  not NOT_50(G88,G89);
  not NOT_51(G90,G91);
  not NOT_52(G92,G93);
  not NOT_53(G94,G95);
  not NOT_54(G96,G95);
  not NOT_55(G97,G98);
  not NOT_56(G99,G88);
  not NOT_57(G17,G94);
  not NOT_58(G100,G101);
  and AND2_0(G102,G103,G16);
  and AND2_1(G104,G16,G82);
  and AND2_2(G105,G20,G82);
  and AND3_0(G106,G24,G22,G82);
  and AND3_1(G107,G62,G18,G82);
  and AND2_3(G108,G95,G51);
  and AND2_4(G3,G81,G90);
  and AND2_5(G109,G110,G51);
  and AND2_6(G1,G80,G92);
  and AND2_7(G111,G96,G110);
  and AND2_8(G112,G96,G113);
  or OR3_0(G114,G20,G18,G16);
  or OR3_1(G115,G24,G22,G60);
  or OR4_0(G116,G62,G22,G20,G16);
  or OR2_0(G117,G65,G60);
  or OR2_1(G118,G72,SPL4_OUT1);
  or OR2_2(G119,G64,G73);
  or OR4_1(G120,G24,G22,G65,G73);
  or OR3_2(G121,G20,G65,G73);
  or OR4_2(G122,G64,G18,G60,G73);
  or OR2_3(G123,G74,SPL1_OUT1);
  or OR4_3(G124,G125,SPL4_OUT2,G18,G64);
  or OR2_4(G87,G126,G34);
  or OR2_5(G127,G128,G36);
  or OR2_6(G129,G76,G38);
  or OR2_7(G130,G79,G43);
  or OR2_8(G131,G83,G42);
  or OR2_9(G98,G132,G26);
  or OR2_10(G133,G134,G28);
  or OR2_11(G135,G136,G30);
  or OR2_12(G137,G84,G32);
  or OR2_13(G101,G138,G18);
  or OR2_14(G139,G140,G20);
  or OR2_15(G141,G142,G22);
  or OR2_16(G143,G99,G24);
  nand NAND2_0(G125,G63,G24);
  nand NAND4_0(G103,G60,G65,G63,G24);
  nand NAND2_1(G144,G128,G36);
  nand NAND2_2(G145,G76,G38);
  nand NAND2_3(G113,G119,G120);
  nand NAND2_4(G146,G121,G122);
  nand NAND2_5(G147,G148,G62);
  nand NAND4_1(G149,G82,G69,G64,G22);
  nand NAND4_2(G150,G82,G20,G117,
    G115);
  nand NAND3_0(G11,G82,G114,G116);
  nand NAND2_6(G151,G152,G124);
  nand NAND2_7(G153,G127,G144);
  nand NAND2_8(G154,G129,G145);
  nand NAND2_9(G91,G130,G118);
  nand NAND3_1(G155,G146,G63,G62);
  nand NAND2_10(G93,G131,G123);
  nand NAND2_11(G95,G151,G147);
  nand NAND2_12(G156,G134,G28);
  nand NAND2_13(G157,G136,G30);
  nand NAND2_14(G158,G84,G32);
  nand NAND2_15(G110,G151,G155);
  nand NAND2_16(G159,G133,G156);
  nand NAND2_17(G160,G135,G157);
  nand NAND2_18(G161,G137,G158);
  nand NAND2_19(G162,G140,G20);
  nand NAND2_20(G163,G142,G22);
  nand NAND2_21(G164,G99,G24);
  nand NAND2_22(G165,G139,G162);
  nand NAND2_23(G166,G141,G163);
  nand NAND2_24(G167,G143,G164);
  nor NOR3_0(G168,G20,G22,G24);
  nor NOR3_1(G169,G36,G38,G40);
  nor NOR3_2(G170,G28,G30,G32);
  nor NOR2_0(G171,G169,G54);
  nor NOR3_3(G126,G55,G56,G57);
  nor NOR2_1(G128,G56,G57);
  nor NOR2_2(G152,G73,G69);
  nor NOR4_0(G148,G73,G60,G64,G22);
  nor NOR2_3(G85,G171,SPL1_OUT2);
  nor NOR3_4(G41,G73,G75,G171);
  nor NOR4_1(G132,G85,G51,G52,G53);
  nor NOR3_5(G134,G85,G52,G53);
  nor NOR3_6(G89,G170,G85,G50);
  nor NOR2_4(G136,G85,G53);
  nor NOR4_2(G13,G104,G105,G106,
    G107);
  nor NOR2_5(G5,G149,G62);
  nor NOR2_6(G15,G150,G102);
  nor NOR3_7(G35,G73,G86,G171);
  nor NOR3_8(G37,G73,G153,G171);
  nor NOR3_9(G39,G73,G154,G171);
  nor NOR4_3(G138,G88,G47,G48,G49);
  nor NOR3_10(G140,G88,G48,G49);
  nor NOR3_11(G172,G168,G88,G46);
  nor NOR2_7(G142,G88,G49);
  nor NOR3_12(G27,G73,G97,G89);
  nor NOR3_13(G29,G73,G159,G89);
  nor NOR3_14(G31,G73,G160,G89);
  nor NOR3_15(G33,G73,G161,G89);
  nor NOR2_8(G9,G111,G109);
  nor NOR2_9(G9,G112,G108);
  nor NOR3_16(G19,G73,G100,G172);
  nor NOR3_17(G21,G73,G165,G172);
  nor NOR3_18(G23,G73,G166,G172);
  nor NOR3_19(G25,G73,G167,G172);

endmodule
